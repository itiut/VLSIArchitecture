module fft064(
              f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
              f_010,f_011,f_012,f_013,f_014,f_015,f_016,f_017,f_018,f_019,
              f_020,f_021,f_022,f_023,f_024,f_025,f_026,f_027,f_028,f_029,
              f_030,f_031,f_032,f_033,f_034,f_035,f_036,f_037,f_038,f_039,
              f_040,f_041,f_042,f_043,f_044,f_045,f_046,f_047,f_048,f_049,
              f_050,f_051,f_052,f_053,f_054,f_055,f_056,f_057,f_058,f_059,
              f_060,f_061,f_062,f_063,
              x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
              x_010,x_011,x_012,x_013,x_014,x_015,x_016,x_017,x_018,x_019,
              x_020,x_021,x_022,x_023,x_024,x_025,x_026,x_027,x_028,x_029,
              x_030,x_031,x_032,x_033,x_034,x_035,x_036,x_037,x_038,x_039,
              x_040,x_041,x_042,x_043,x_044,x_045,x_046,x_047,x_048,x_049,
              x_050,x_051,x_052,x_053,x_054,x_055,x_056,x_057,x_058,x_059,
              x_060,x_061,x_062,x_063,
              W000,W001,W002,W003,W004,W005,W006,W007,W008,W009,
              W010,W011,W012,W013,W014,W015,W016,W017,W018,W019,
              W020,W021,W022,W023,W024,W025,W026,W027,W028,W029,
              W030,W031);
    output [31:0]
                  f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
                  f_010,f_011,f_012,f_013,f_014,f_015,f_016,f_017,f_018,f_019,
                  f_020,f_021,f_022,f_023,f_024,f_025,f_026,f_027,f_028,f_029,
                  f_030,f_031,f_032,f_033,f_034,f_035,f_036,f_037,f_038,f_039,
                  f_040,f_041,f_042,f_043,f_044,f_045,f_046,f_047,f_048,f_049,
                  f_050,f_051,f_052,f_053,f_054,f_055,f_056,f_057,f_058,f_059,
                  f_060,f_061,f_062,f_063;
    input [31:0]
                 x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
                 x_010,x_011,x_012,x_013,x_014,x_015,x_016,x_017,x_018,x_019,
                 x_020,x_021,x_022,x_023,x_024,x_025,x_026,x_027,x_028,x_029,
                 x_030,x_031,x_032,x_033,x_034,x_035,x_036,x_037,x_038,x_039,
                 x_040,x_041,x_042,x_043,x_044,x_045,x_046,x_047,x_048,x_049,
                 x_050,x_051,x_052,x_053,x_054,x_055,x_056,x_057,x_058,x_059,
                 x_060,x_061,x_062,x_063;
    input [31:0]
                 W000,W001,W002,W003,W004,W005,W006,W007,W008,W009,
                 W010,W011,W012,W013,W014,W015,W016,W017,W018,W019,
                 W020,W021,W022,W023,W024,W025,W026,W027,W028,W029,
                 W030,W031;
    wire [31:0]
               x_00_000,x_00_001,x_00_002,x_00_003,x_00_004,x_00_005,x_00_006,x_00_007,x_00_008,x_00_009,
               x_00_010,x_00_011,x_00_012,x_00_013,x_00_014,x_00_015,x_00_016,x_00_017,x_00_018,x_00_019,
               x_00_020,x_00_021,x_00_022,x_00_023,x_00_024,x_00_025,x_00_026,x_00_027,x_00_028,x_00_029,
               x_00_030,x_00_031,x_00_032,x_00_033,x_00_034,x_00_035,x_00_036,x_00_037,x_00_038,x_00_039,
               x_00_040,x_00_041,x_00_042,x_00_043,x_00_044,x_00_045,x_00_046,x_00_047,x_00_048,x_00_049,
               x_00_050,x_00_051,x_00_052,x_00_053,x_00_054,x_00_055,x_00_056,x_00_057,x_00_058,x_00_059,
               x_00_060,x_00_061,x_00_062,x_00_063,
               x_01_000,x_01_001,x_01_002,x_01_003,x_01_004,x_01_005,x_01_006,x_01_007,x_01_008,x_01_009,
               x_01_010,x_01_011,x_01_012,x_01_013,x_01_014,x_01_015,x_01_016,x_01_017,x_01_018,x_01_019,
               x_01_020,x_01_021,x_01_022,x_01_023,x_01_024,x_01_025,x_01_026,x_01_027,x_01_028,x_01_029,
               x_01_030,x_01_031,x_01_032,x_01_033,x_01_034,x_01_035,x_01_036,x_01_037,x_01_038,x_01_039,
               x_01_040,x_01_041,x_01_042,x_01_043,x_01_044,x_01_045,x_01_046,x_01_047,x_01_048,x_01_049,
               x_01_050,x_01_051,x_01_052,x_01_053,x_01_054,x_01_055,x_01_056,x_01_057,x_01_058,x_01_059,
               x_01_060,x_01_061,x_01_062,x_01_063,
               x_02_000,x_02_001,x_02_002,x_02_003,x_02_004,x_02_005,x_02_006,x_02_007,x_02_008,x_02_009,
               x_02_010,x_02_011,x_02_012,x_02_013,x_02_014,x_02_015,x_02_016,x_02_017,x_02_018,x_02_019,
               x_02_020,x_02_021,x_02_022,x_02_023,x_02_024,x_02_025,x_02_026,x_02_027,x_02_028,x_02_029,
               x_02_030,x_02_031,x_02_032,x_02_033,x_02_034,x_02_035,x_02_036,x_02_037,x_02_038,x_02_039,
               x_02_040,x_02_041,x_02_042,x_02_043,x_02_044,x_02_045,x_02_046,x_02_047,x_02_048,x_02_049,
               x_02_050,x_02_051,x_02_052,x_02_053,x_02_054,x_02_055,x_02_056,x_02_057,x_02_058,x_02_059,
               x_02_060,x_02_061,x_02_062,x_02_063,
               x_03_000,x_03_001,x_03_002,x_03_003,x_03_004,x_03_005,x_03_006,x_03_007,x_03_008,x_03_009,
               x_03_010,x_03_011,x_03_012,x_03_013,x_03_014,x_03_015,x_03_016,x_03_017,x_03_018,x_03_019,
               x_03_020,x_03_021,x_03_022,x_03_023,x_03_024,x_03_025,x_03_026,x_03_027,x_03_028,x_03_029,
               x_03_030,x_03_031,x_03_032,x_03_033,x_03_034,x_03_035,x_03_036,x_03_037,x_03_038,x_03_039,
               x_03_040,x_03_041,x_03_042,x_03_043,x_03_044,x_03_045,x_03_046,x_03_047,x_03_048,x_03_049,
               x_03_050,x_03_051,x_03_052,x_03_053,x_03_054,x_03_055,x_03_056,x_03_057,x_03_058,x_03_059,
               x_03_060,x_03_061,x_03_062,x_03_063,
               x_04_000,x_04_001,x_04_002,x_04_003,x_04_004,x_04_005,x_04_006,x_04_007,x_04_008,x_04_009,
               x_04_010,x_04_011,x_04_012,x_04_013,x_04_014,x_04_015,x_04_016,x_04_017,x_04_018,x_04_019,
               x_04_020,x_04_021,x_04_022,x_04_023,x_04_024,x_04_025,x_04_026,x_04_027,x_04_028,x_04_029,
               x_04_030,x_04_031,x_04_032,x_04_033,x_04_034,x_04_035,x_04_036,x_04_037,x_04_038,x_04_039,
               x_04_040,x_04_041,x_04_042,x_04_043,x_04_044,x_04_045,x_04_046,x_04_047,x_04_048,x_04_049,
               x_04_050,x_04_051,x_04_052,x_04_053,x_04_054,x_04_055,x_04_056,x_04_057,x_04_058,x_04_059,
               x_04_060,x_04_061,x_04_062,x_04_063,
               x_05_000,x_05_001,x_05_002,x_05_003,x_05_004,x_05_005,x_05_006,x_05_007,x_05_008,x_05_009,
               x_05_010,x_05_011,x_05_012,x_05_013,x_05_014,x_05_015,x_05_016,x_05_017,x_05_018,x_05_019,
               x_05_020,x_05_021,x_05_022,x_05_023,x_05_024,x_05_025,x_05_026,x_05_027,x_05_028,x_05_029,
               x_05_030,x_05_031,x_05_032,x_05_033,x_05_034,x_05_035,x_05_036,x_05_037,x_05_038,x_05_039,
               x_05_040,x_05_041,x_05_042,x_05_043,x_05_044,x_05_045,x_05_046,x_05_047,x_05_048,x_05_049,
               x_05_050,x_05_051,x_05_052,x_05_053,x_05_054,x_05_055,x_05_056,x_05_057,x_05_058,x_05_059,
               x_05_060,x_05_061,x_05_062,x_05_063,
               x_06_000,x_06_001,x_06_002,x_06_003,x_06_004,x_06_005,x_06_006,x_06_007,x_06_008,x_06_009,
               x_06_010,x_06_011,x_06_012,x_06_013,x_06_014,x_06_015,x_06_016,x_06_017,x_06_018,x_06_019,
               x_06_020,x_06_021,x_06_022,x_06_023,x_06_024,x_06_025,x_06_026,x_06_027,x_06_028,x_06_029,
               x_06_030,x_06_031,x_06_032,x_06_033,x_06_034,x_06_035,x_06_036,x_06_037,x_06_038,x_06_039,
               x_06_040,x_06_041,x_06_042,x_06_043,x_06_044,x_06_045,x_06_046,x_06_047,x_06_048,x_06_049,
               x_06_050,x_06_051,x_06_052,x_06_053,x_06_054,x_06_055,x_06_056,x_06_057,x_06_058,x_06_059,
               x_06_060,x_06_061,x_06_062,x_06_063;
    assign x_00_000 = x_000;
    assign x_00_001 = x_001;
    assign x_00_002 = x_002;
    assign x_00_003 = x_003;
    assign x_00_004 = x_004;
    assign x_00_005 = x_005;
    assign x_00_006 = x_006;
    assign x_00_007 = x_007;
    assign x_00_008 = x_008;
    assign x_00_009 = x_009;
    assign x_00_010 = x_010;
    assign x_00_011 = x_011;
    assign x_00_012 = x_012;
    assign x_00_013 = x_013;
    assign x_00_014 = x_014;
    assign x_00_015 = x_015;
    assign x_00_016 = x_016;
    assign x_00_017 = x_017;
    assign x_00_018 = x_018;
    assign x_00_019 = x_019;
    assign x_00_020 = x_020;
    assign x_00_021 = x_021;
    assign x_00_022 = x_022;
    assign x_00_023 = x_023;
    assign x_00_024 = x_024;
    assign x_00_025 = x_025;
    assign x_00_026 = x_026;
    assign x_00_027 = x_027;
    assign x_00_028 = x_028;
    assign x_00_029 = x_029;
    assign x_00_030 = x_030;
    assign x_00_031 = x_031;
    assign x_00_032 = x_032;
    assign x_00_033 = x_033;
    assign x_00_034 = x_034;
    assign x_00_035 = x_035;
    assign x_00_036 = x_036;
    assign x_00_037 = x_037;
    assign x_00_038 = x_038;
    assign x_00_039 = x_039;
    assign x_00_040 = x_040;
    assign x_00_041 = x_041;
    assign x_00_042 = x_042;
    assign x_00_043 = x_043;
    assign x_00_044 = x_044;
    assign x_00_045 = x_045;
    assign x_00_046 = x_046;
    assign x_00_047 = x_047;
    assign x_00_048 = x_048;
    assign x_00_049 = x_049;
    assign x_00_050 = x_050;
    assign x_00_051 = x_051;
    assign x_00_052 = x_052;
    assign x_00_053 = x_053;
    assign x_00_054 = x_054;
    assign x_00_055 = x_055;
    assign x_00_056 = x_056;
    assign x_00_057 = x_057;
    assign x_00_058 = x_058;
    assign x_00_059 = x_059;
    assign x_00_060 = x_060;
    assign x_00_061 = x_061;
    assign x_00_062 = x_062;
    assign x_00_063 = x_063;
    assign x_00_000 = x_000;
    assign x_00_001 = x_001;
    assign x_00_002 = x_002;
    assign x_00_003 = x_003;
    assign x_00_004 = x_004;
    assign x_00_005 = x_005;
    assign x_00_006 = x_006;
    assign x_00_007 = x_007;
    assign x_00_008 = x_008;
    assign x_00_009 = x_009;
    assign x_00_010 = x_010;
    assign x_00_011 = x_011;
    assign x_00_012 = x_012;
    assign x_00_013 = x_013;
    assign x_00_014 = x_014;
    assign x_00_015 = x_015;
    assign x_00_016 = x_016;
    assign x_00_017 = x_017;
    assign x_00_018 = x_018;
    assign x_00_019 = x_019;
    assign x_00_020 = x_020;
    assign x_00_021 = x_021;
    assign x_00_022 = x_022;
    assign x_00_023 = x_023;
    assign x_00_024 = x_024;
    assign x_00_025 = x_025;
    assign x_00_026 = x_026;
    assign x_00_027 = x_027;
    assign x_00_028 = x_028;
    assign x_00_029 = x_029;
    assign x_00_030 = x_030;
    assign x_00_031 = x_031;
    assign x_00_032 = x_032;
    assign x_00_033 = x_033;
    assign x_00_034 = x_034;
    assign x_00_035 = x_035;
    assign x_00_036 = x_036;
    assign x_00_037 = x_037;
    assign x_00_038 = x_038;
    assign x_00_039 = x_039;
    assign x_00_040 = x_040;
    assign x_00_041 = x_041;
    assign x_00_042 = x_042;
    assign x_00_043 = x_043;
    assign x_00_044 = x_044;
    assign x_00_045 = x_045;
    assign x_00_046 = x_046;
    assign x_00_047 = x_047;
    assign x_00_048 = x_048;
    assign x_00_049 = x_049;
    assign x_00_050 = x_050;
    assign x_00_051 = x_051;
    assign x_00_052 = x_052;
    assign x_00_053 = x_053;
    assign x_00_054 = x_054;
    assign x_00_055 = x_055;
    assign x_00_056 = x_056;
    assign x_00_057 = x_057;
    assign x_00_058 = x_058;
    assign x_00_059 = x_059;
    assign x_00_060 = x_060;
    assign x_00_061 = x_061;
    assign x_00_062 = x_062;
    assign x_00_063 = x_063;
    butt2 xx_00_000( .x0(x_00_000), .x1(x_00_032), .y0(x_01_000), .y1(x_01_032), .W(W000) );
    butt2 xx_00_001( .x0(x_00_016), .x1(x_00_048), .y0(x_01_016), .y1(x_01_048), .W(W000) );
    butt2 xx_00_002( .x0(x_00_008), .x1(x_00_040), .y0(x_01_008), .y1(x_01_040), .W(W000) );
    butt2 xx_00_003( .x0(x_00_024), .x1(x_00_056), .y0(x_01_024), .y1(x_01_056), .W(W000) );
    butt2 xx_00_004( .x0(x_00_004), .x1(x_00_036), .y0(x_01_004), .y1(x_01_036), .W(W000) );
    butt2 xx_00_005( .x0(x_00_020), .x1(x_00_052), .y0(x_01_020), .y1(x_01_052), .W(W000) );
    butt2 xx_00_006( .x0(x_00_012), .x1(x_00_044), .y0(x_01_012), .y1(x_01_044), .W(W000) );
    butt2 xx_00_007( .x0(x_00_028), .x1(x_00_060), .y0(x_01_028), .y1(x_01_060), .W(W000) );
    butt2 xx_00_008( .x0(x_00_002), .x1(x_00_034), .y0(x_01_002), .y1(x_01_034), .W(W000) );
    butt2 xx_00_009( .x0(x_00_018), .x1(x_00_050), .y0(x_01_018), .y1(x_01_050), .W(W000) );
    butt2 xx_00_010( .x0(x_00_010), .x1(x_00_042), .y0(x_01_010), .y1(x_01_042), .W(W000) );
    butt2 xx_00_011( .x0(x_00_026), .x1(x_00_058), .y0(x_01_026), .y1(x_01_058), .W(W000) );
    butt2 xx_00_012( .x0(x_00_006), .x1(x_00_038), .y0(x_01_006), .y1(x_01_038), .W(W000) );
    butt2 xx_00_013( .x0(x_00_022), .x1(x_00_054), .y0(x_01_022), .y1(x_01_054), .W(W000) );
    butt2 xx_00_014( .x0(x_00_014), .x1(x_00_046), .y0(x_01_014), .y1(x_01_046), .W(W000) );
    butt2 xx_00_015( .x0(x_00_030), .x1(x_00_062), .y0(x_01_030), .y1(x_01_062), .W(W000) );
    butt2 xx_00_016( .x0(x_00_001), .x1(x_00_033), .y0(x_01_001), .y1(x_01_033), .W(W000) );
    butt2 xx_00_017( .x0(x_00_017), .x1(x_00_049), .y0(x_01_017), .y1(x_01_049), .W(W000) );
    butt2 xx_00_018( .x0(x_00_009), .x1(x_00_041), .y0(x_01_009), .y1(x_01_041), .W(W000) );
    butt2 xx_00_019( .x0(x_00_025), .x1(x_00_057), .y0(x_01_025), .y1(x_01_057), .W(W000) );
    butt2 xx_00_020( .x0(x_00_005), .x1(x_00_037), .y0(x_01_005), .y1(x_01_037), .W(W000) );
    butt2 xx_00_021( .x0(x_00_021), .x1(x_00_053), .y0(x_01_021), .y1(x_01_053), .W(W000) );
    butt2 xx_00_022( .x0(x_00_013), .x1(x_00_045), .y0(x_01_013), .y1(x_01_045), .W(W000) );
    butt2 xx_00_023( .x0(x_00_029), .x1(x_00_061), .y0(x_01_029), .y1(x_01_061), .W(W000) );
    butt2 xx_00_024( .x0(x_00_003), .x1(x_00_035), .y0(x_01_003), .y1(x_01_035), .W(W000) );
    butt2 xx_00_025( .x0(x_00_019), .x1(x_00_051), .y0(x_01_019), .y1(x_01_051), .W(W000) );
    butt2 xx_00_026( .x0(x_00_011), .x1(x_00_043), .y0(x_01_011), .y1(x_01_043), .W(W000) );
    butt2 xx_00_027( .x0(x_00_027), .x1(x_00_059), .y0(x_01_027), .y1(x_01_059), .W(W000) );
    butt2 xx_00_028( .x0(x_00_007), .x1(x_00_039), .y0(x_01_007), .y1(x_01_039), .W(W000) );
    butt2 xx_00_029( .x0(x_00_023), .x1(x_00_055), .y0(x_01_023), .y1(x_01_055), .W(W000) );
    butt2 xx_00_030( .x0(x_00_015), .x1(x_00_047), .y0(x_01_015), .y1(x_01_047), .W(W000) );
    butt2 xx_00_031( .x0(x_00_031), .x1(x_00_063), .y0(x_01_031), .y1(x_01_063), .W(W000) );
    butt2 xx_01_000( .x0(x_01_000), .x1(x_01_016), .y0(x_02_000), .y1(x_02_016), .W(W000) );
    butt2 xx_01_001( .x0(x_01_032), .x1(x_01_048), .y0(x_02_032), .y1(x_02_048), .W(W016) );
    butt2 xx_01_002( .x0(x_01_008), .x1(x_01_024), .y0(x_02_008), .y1(x_02_024), .W(W000) );
    butt2 xx_01_003( .x0(x_01_040), .x1(x_01_056), .y0(x_02_040), .y1(x_02_056), .W(W016) );
    butt2 xx_01_004( .x0(x_01_004), .x1(x_01_020), .y0(x_02_004), .y1(x_02_020), .W(W000) );
    butt2 xx_01_005( .x0(x_01_036), .x1(x_01_052), .y0(x_02_036), .y1(x_02_052), .W(W016) );
    butt2 xx_01_006( .x0(x_01_012), .x1(x_01_028), .y0(x_02_012), .y1(x_02_028), .W(W000) );
    butt2 xx_01_007( .x0(x_01_044), .x1(x_01_060), .y0(x_02_044), .y1(x_02_060), .W(W016) );
    butt2 xx_01_008( .x0(x_01_002), .x1(x_01_018), .y0(x_02_002), .y1(x_02_018), .W(W000) );
    butt2 xx_01_009( .x0(x_01_034), .x1(x_01_050), .y0(x_02_034), .y1(x_02_050), .W(W016) );
    butt2 xx_01_010( .x0(x_01_010), .x1(x_01_026), .y0(x_02_010), .y1(x_02_026), .W(W000) );
    butt2 xx_01_011( .x0(x_01_042), .x1(x_01_058), .y0(x_02_042), .y1(x_02_058), .W(W016) );
    butt2 xx_01_012( .x0(x_01_006), .x1(x_01_022), .y0(x_02_006), .y1(x_02_022), .W(W000) );
    butt2 xx_01_013( .x0(x_01_038), .x1(x_01_054), .y0(x_02_038), .y1(x_02_054), .W(W016) );
    butt2 xx_01_014( .x0(x_01_014), .x1(x_01_030), .y0(x_02_014), .y1(x_02_030), .W(W000) );
    butt2 xx_01_015( .x0(x_01_046), .x1(x_01_062), .y0(x_02_046), .y1(x_02_062), .W(W016) );
    butt2 xx_01_016( .x0(x_01_001), .x1(x_01_017), .y0(x_02_001), .y1(x_02_017), .W(W000) );
    butt2 xx_01_017( .x0(x_01_033), .x1(x_01_049), .y0(x_02_033), .y1(x_02_049), .W(W016) );
    butt2 xx_01_018( .x0(x_01_009), .x1(x_01_025), .y0(x_02_009), .y1(x_02_025), .W(W000) );
    butt2 xx_01_019( .x0(x_01_041), .x1(x_01_057), .y0(x_02_041), .y1(x_02_057), .W(W016) );
    butt2 xx_01_020( .x0(x_01_005), .x1(x_01_021), .y0(x_02_005), .y1(x_02_021), .W(W000) );
    butt2 xx_01_021( .x0(x_01_037), .x1(x_01_053), .y0(x_02_037), .y1(x_02_053), .W(W016) );
    butt2 xx_01_022( .x0(x_01_013), .x1(x_01_029), .y0(x_02_013), .y1(x_02_029), .W(W000) );
    butt2 xx_01_023( .x0(x_01_045), .x1(x_01_061), .y0(x_02_045), .y1(x_02_061), .W(W016) );
    butt2 xx_01_024( .x0(x_01_003), .x1(x_01_019), .y0(x_02_003), .y1(x_02_019), .W(W000) );
    butt2 xx_01_025( .x0(x_01_035), .x1(x_01_051), .y0(x_02_035), .y1(x_02_051), .W(W016) );
    butt2 xx_01_026( .x0(x_01_011), .x1(x_01_027), .y0(x_02_011), .y1(x_02_027), .W(W000) );
    butt2 xx_01_027( .x0(x_01_043), .x1(x_01_059), .y0(x_02_043), .y1(x_02_059), .W(W016) );
    butt2 xx_01_028( .x0(x_01_007), .x1(x_01_023), .y0(x_02_007), .y1(x_02_023), .W(W000) );
    butt2 xx_01_029( .x0(x_01_039), .x1(x_01_055), .y0(x_02_039), .y1(x_02_055), .W(W016) );
    butt2 xx_01_030( .x0(x_01_015), .x1(x_01_031), .y0(x_02_015), .y1(x_02_031), .W(W000) );
    butt2 xx_01_031( .x0(x_01_047), .x1(x_01_063), .y0(x_02_047), .y1(x_02_063), .W(W016) );
    butt2 xx_02_000( .x0(x_02_000), .x1(x_02_008), .y0(x_03_000), .y1(x_03_008), .W(W000) );
    butt2 xx_02_001( .x0(x_02_032), .x1(x_02_040), .y0(x_03_032), .y1(x_03_040), .W(W008) );
    butt2 xx_02_002( .x0(x_02_016), .x1(x_02_024), .y0(x_03_016), .y1(x_03_024), .W(W016) );
    butt2 xx_02_003( .x0(x_02_048), .x1(x_02_056), .y0(x_03_048), .y1(x_03_056), .W(W024) );
    butt2 xx_02_004( .x0(x_02_004), .x1(x_02_012), .y0(x_03_004), .y1(x_03_012), .W(W000) );
    butt2 xx_02_005( .x0(x_02_036), .x1(x_02_044), .y0(x_03_036), .y1(x_03_044), .W(W008) );
    butt2 xx_02_006( .x0(x_02_020), .x1(x_02_028), .y0(x_03_020), .y1(x_03_028), .W(W016) );
    butt2 xx_02_007( .x0(x_02_052), .x1(x_02_060), .y0(x_03_052), .y1(x_03_060), .W(W024) );
    butt2 xx_02_008( .x0(x_02_002), .x1(x_02_010), .y0(x_03_002), .y1(x_03_010), .W(W000) );
    butt2 xx_02_009( .x0(x_02_034), .x1(x_02_042), .y0(x_03_034), .y1(x_03_042), .W(W008) );
    butt2 xx_02_010( .x0(x_02_018), .x1(x_02_026), .y0(x_03_018), .y1(x_03_026), .W(W016) );
    butt2 xx_02_011( .x0(x_02_050), .x1(x_02_058), .y0(x_03_050), .y1(x_03_058), .W(W024) );
    butt2 xx_02_012( .x0(x_02_006), .x1(x_02_014), .y0(x_03_006), .y1(x_03_014), .W(W000) );
    butt2 xx_02_013( .x0(x_02_038), .x1(x_02_046), .y0(x_03_038), .y1(x_03_046), .W(W008) );
    butt2 xx_02_014( .x0(x_02_022), .x1(x_02_030), .y0(x_03_022), .y1(x_03_030), .W(W016) );
    butt2 xx_02_015( .x0(x_02_054), .x1(x_02_062), .y0(x_03_054), .y1(x_03_062), .W(W024) );
    butt2 xx_02_016( .x0(x_02_001), .x1(x_02_009), .y0(x_03_001), .y1(x_03_009), .W(W000) );
    butt2 xx_02_017( .x0(x_02_033), .x1(x_02_041), .y0(x_03_033), .y1(x_03_041), .W(W008) );
    butt2 xx_02_018( .x0(x_02_017), .x1(x_02_025), .y0(x_03_017), .y1(x_03_025), .W(W016) );
    butt2 xx_02_019( .x0(x_02_049), .x1(x_02_057), .y0(x_03_049), .y1(x_03_057), .W(W024) );
    butt2 xx_02_020( .x0(x_02_005), .x1(x_02_013), .y0(x_03_005), .y1(x_03_013), .W(W000) );
    butt2 xx_02_021( .x0(x_02_037), .x1(x_02_045), .y0(x_03_037), .y1(x_03_045), .W(W008) );
    butt2 xx_02_022( .x0(x_02_021), .x1(x_02_029), .y0(x_03_021), .y1(x_03_029), .W(W016) );
    butt2 xx_02_023( .x0(x_02_053), .x1(x_02_061), .y0(x_03_053), .y1(x_03_061), .W(W024) );
    butt2 xx_02_024( .x0(x_02_003), .x1(x_02_011), .y0(x_03_003), .y1(x_03_011), .W(W000) );
    butt2 xx_02_025( .x0(x_02_035), .x1(x_02_043), .y0(x_03_035), .y1(x_03_043), .W(W008) );
    butt2 xx_02_026( .x0(x_02_019), .x1(x_02_027), .y0(x_03_019), .y1(x_03_027), .W(W016) );
    butt2 xx_02_027( .x0(x_02_051), .x1(x_02_059), .y0(x_03_051), .y1(x_03_059), .W(W024) );
    butt2 xx_02_028( .x0(x_02_007), .x1(x_02_015), .y0(x_03_007), .y1(x_03_015), .W(W000) );
    butt2 xx_02_029( .x0(x_02_039), .x1(x_02_047), .y0(x_03_039), .y1(x_03_047), .W(W008) );
    butt2 xx_02_030( .x0(x_02_023), .x1(x_02_031), .y0(x_03_023), .y1(x_03_031), .W(W016) );
    butt2 xx_02_031( .x0(x_02_055), .x1(x_02_063), .y0(x_03_055), .y1(x_03_063), .W(W024) );
    butt2 xx_03_000( .x0(x_03_000), .x1(x_03_004), .y0(x_04_000), .y1(x_04_004), .W(W000) );
    butt2 xx_03_001( .x0(x_03_032), .x1(x_03_036), .y0(x_04_032), .y1(x_04_036), .W(W004) );
    butt2 xx_03_002( .x0(x_03_016), .x1(x_03_020), .y0(x_04_016), .y1(x_04_020), .W(W008) );
    butt2 xx_03_003( .x0(x_03_048), .x1(x_03_052), .y0(x_04_048), .y1(x_04_052), .W(W012) );
    butt2 xx_03_004( .x0(x_03_008), .x1(x_03_012), .y0(x_04_008), .y1(x_04_012), .W(W016) );
    butt2 xx_03_005( .x0(x_03_040), .x1(x_03_044), .y0(x_04_040), .y1(x_04_044), .W(W020) );
    butt2 xx_03_006( .x0(x_03_024), .x1(x_03_028), .y0(x_04_024), .y1(x_04_028), .W(W024) );
    butt2 xx_03_007( .x0(x_03_056), .x1(x_03_060), .y0(x_04_056), .y1(x_04_060), .W(W028) );
    butt2 xx_03_008( .x0(x_03_002), .x1(x_03_006), .y0(x_04_002), .y1(x_04_006), .W(W000) );
    butt2 xx_03_009( .x0(x_03_034), .x1(x_03_038), .y0(x_04_034), .y1(x_04_038), .W(W004) );
    butt2 xx_03_010( .x0(x_03_018), .x1(x_03_022), .y0(x_04_018), .y1(x_04_022), .W(W008) );
    butt2 xx_03_011( .x0(x_03_050), .x1(x_03_054), .y0(x_04_050), .y1(x_04_054), .W(W012) );
    butt2 xx_03_012( .x0(x_03_010), .x1(x_03_014), .y0(x_04_010), .y1(x_04_014), .W(W016) );
    butt2 xx_03_013( .x0(x_03_042), .x1(x_03_046), .y0(x_04_042), .y1(x_04_046), .W(W020) );
    butt2 xx_03_014( .x0(x_03_026), .x1(x_03_030), .y0(x_04_026), .y1(x_04_030), .W(W024) );
    butt2 xx_03_015( .x0(x_03_058), .x1(x_03_062), .y0(x_04_058), .y1(x_04_062), .W(W028) );
    butt2 xx_03_016( .x0(x_03_001), .x1(x_03_005), .y0(x_04_001), .y1(x_04_005), .W(W000) );
    butt2 xx_03_017( .x0(x_03_033), .x1(x_03_037), .y0(x_04_033), .y1(x_04_037), .W(W004) );
    butt2 xx_03_018( .x0(x_03_017), .x1(x_03_021), .y0(x_04_017), .y1(x_04_021), .W(W008) );
    butt2 xx_03_019( .x0(x_03_049), .x1(x_03_053), .y0(x_04_049), .y1(x_04_053), .W(W012) );
    butt2 xx_03_020( .x0(x_03_009), .x1(x_03_013), .y0(x_04_009), .y1(x_04_013), .W(W016) );
    butt2 xx_03_021( .x0(x_03_041), .x1(x_03_045), .y0(x_04_041), .y1(x_04_045), .W(W020) );
    butt2 xx_03_022( .x0(x_03_025), .x1(x_03_029), .y0(x_04_025), .y1(x_04_029), .W(W024) );
    butt2 xx_03_023( .x0(x_03_057), .x1(x_03_061), .y0(x_04_057), .y1(x_04_061), .W(W028) );
    butt2 xx_03_024( .x0(x_03_003), .x1(x_03_007), .y0(x_04_003), .y1(x_04_007), .W(W000) );
    butt2 xx_03_025( .x0(x_03_035), .x1(x_03_039), .y0(x_04_035), .y1(x_04_039), .W(W004) );
    butt2 xx_03_026( .x0(x_03_019), .x1(x_03_023), .y0(x_04_019), .y1(x_04_023), .W(W008) );
    butt2 xx_03_027( .x0(x_03_051), .x1(x_03_055), .y0(x_04_051), .y1(x_04_055), .W(W012) );
    butt2 xx_03_028( .x0(x_03_011), .x1(x_03_015), .y0(x_04_011), .y1(x_04_015), .W(W016) );
    butt2 xx_03_029( .x0(x_03_043), .x1(x_03_047), .y0(x_04_043), .y1(x_04_047), .W(W020) );
    butt2 xx_03_030( .x0(x_03_027), .x1(x_03_031), .y0(x_04_027), .y1(x_04_031), .W(W024) );
    butt2 xx_03_031( .x0(x_03_059), .x1(x_03_063), .y0(x_04_059), .y1(x_04_063), .W(W028) );
    butt2 xx_04_000( .x0(x_04_000), .x1(x_04_002), .y0(x_05_000), .y1(x_05_002), .W(W000) );
    butt2 xx_04_001( .x0(x_04_032), .x1(x_04_034), .y0(x_05_032), .y1(x_05_034), .W(W002) );
    butt2 xx_04_002( .x0(x_04_016), .x1(x_04_018), .y0(x_05_016), .y1(x_05_018), .W(W004) );
    butt2 xx_04_003( .x0(x_04_048), .x1(x_04_050), .y0(x_05_048), .y1(x_05_050), .W(W006) );
    butt2 xx_04_004( .x0(x_04_008), .x1(x_04_010), .y0(x_05_008), .y1(x_05_010), .W(W008) );
    butt2 xx_04_005( .x0(x_04_040), .x1(x_04_042), .y0(x_05_040), .y1(x_05_042), .W(W010) );
    butt2 xx_04_006( .x0(x_04_024), .x1(x_04_026), .y0(x_05_024), .y1(x_05_026), .W(W012) );
    butt2 xx_04_007( .x0(x_04_056), .x1(x_04_058), .y0(x_05_056), .y1(x_05_058), .W(W014) );
    butt2 xx_04_008( .x0(x_04_004), .x1(x_04_006), .y0(x_05_004), .y1(x_05_006), .W(W016) );
    butt2 xx_04_009( .x0(x_04_036), .x1(x_04_038), .y0(x_05_036), .y1(x_05_038), .W(W018) );
    butt2 xx_04_010( .x0(x_04_020), .x1(x_04_022), .y0(x_05_020), .y1(x_05_022), .W(W020) );
    butt2 xx_04_011( .x0(x_04_052), .x1(x_04_054), .y0(x_05_052), .y1(x_05_054), .W(W022) );
    butt2 xx_04_012( .x0(x_04_012), .x1(x_04_014), .y0(x_05_012), .y1(x_05_014), .W(W024) );
    butt2 xx_04_013( .x0(x_04_044), .x1(x_04_046), .y0(x_05_044), .y1(x_05_046), .W(W026) );
    butt2 xx_04_014( .x0(x_04_028), .x1(x_04_030), .y0(x_05_028), .y1(x_05_030), .W(W028) );
    butt2 xx_04_015( .x0(x_04_060), .x1(x_04_062), .y0(x_05_060), .y1(x_05_062), .W(W030) );
    butt2 xx_04_016( .x0(x_04_001), .x1(x_04_003), .y0(x_05_001), .y1(x_05_003), .W(W000) );
    butt2 xx_04_017( .x0(x_04_033), .x1(x_04_035), .y0(x_05_033), .y1(x_05_035), .W(W002) );
    butt2 xx_04_018( .x0(x_04_017), .x1(x_04_019), .y0(x_05_017), .y1(x_05_019), .W(W004) );
    butt2 xx_04_019( .x0(x_04_049), .x1(x_04_051), .y0(x_05_049), .y1(x_05_051), .W(W006) );
    butt2 xx_04_020( .x0(x_04_009), .x1(x_04_011), .y0(x_05_009), .y1(x_05_011), .W(W008) );
    butt2 xx_04_021( .x0(x_04_041), .x1(x_04_043), .y0(x_05_041), .y1(x_05_043), .W(W010) );
    butt2 xx_04_022( .x0(x_04_025), .x1(x_04_027), .y0(x_05_025), .y1(x_05_027), .W(W012) );
    butt2 xx_04_023( .x0(x_04_057), .x1(x_04_059), .y0(x_05_057), .y1(x_05_059), .W(W014) );
    butt2 xx_04_024( .x0(x_04_005), .x1(x_04_007), .y0(x_05_005), .y1(x_05_007), .W(W016) );
    butt2 xx_04_025( .x0(x_04_037), .x1(x_04_039), .y0(x_05_037), .y1(x_05_039), .W(W018) );
    butt2 xx_04_026( .x0(x_04_021), .x1(x_04_023), .y0(x_05_021), .y1(x_05_023), .W(W020) );
    butt2 xx_04_027( .x0(x_04_053), .x1(x_04_055), .y0(x_05_053), .y1(x_05_055), .W(W022) );
    butt2 xx_04_028( .x0(x_04_013), .x1(x_04_015), .y0(x_05_013), .y1(x_05_015), .W(W024) );
    butt2 xx_04_029( .x0(x_04_045), .x1(x_04_047), .y0(x_05_045), .y1(x_05_047), .W(W026) );
    butt2 xx_04_030( .x0(x_04_029), .x1(x_04_031), .y0(x_05_029), .y1(x_05_031), .W(W028) );
    butt2 xx_04_031( .x0(x_04_061), .x1(x_04_063), .y0(x_05_061), .y1(x_05_063), .W(W030) );
    butt2 xx_05_000( .x0(x_05_000), .x1(x_05_001), .y0(x_06_000), .y1(x_06_001), .W(W000) );
    assign f_000 = x_06_000;
    assign f_032 = x_06_001;
    butt2 xx_05_001( .x0(x_05_032), .x1(x_05_033), .y0(x_06_032), .y1(x_06_033), .W(W001) );
    assign f_001 = x_06_032;
    assign f_033 = x_06_033;
    butt2 xx_05_002( .x0(x_05_016), .x1(x_05_017), .y0(x_06_016), .y1(x_06_017), .W(W002) );
    assign f_002 = x_06_016;
    assign f_034 = x_06_017;
    butt2 xx_05_003( .x0(x_05_048), .x1(x_05_049), .y0(x_06_048), .y1(x_06_049), .W(W003) );
    assign f_003 = x_06_048;
    assign f_035 = x_06_049;
    butt2 xx_05_004( .x0(x_05_008), .x1(x_05_009), .y0(x_06_008), .y1(x_06_009), .W(W004) );
    assign f_004 = x_06_008;
    assign f_036 = x_06_009;
    butt2 xx_05_005( .x0(x_05_040), .x1(x_05_041), .y0(x_06_040), .y1(x_06_041), .W(W005) );
    assign f_005 = x_06_040;
    assign f_037 = x_06_041;
    butt2 xx_05_006( .x0(x_05_024), .x1(x_05_025), .y0(x_06_024), .y1(x_06_025), .W(W006) );
    assign f_006 = x_06_024;
    assign f_038 = x_06_025;
    butt2 xx_05_007( .x0(x_05_056), .x1(x_05_057), .y0(x_06_056), .y1(x_06_057), .W(W007) );
    assign f_007 = x_06_056;
    assign f_039 = x_06_057;
    butt2 xx_05_008( .x0(x_05_004), .x1(x_05_005), .y0(x_06_004), .y1(x_06_005), .W(W008) );
    assign f_008 = x_06_004;
    assign f_040 = x_06_005;
    butt2 xx_05_009( .x0(x_05_036), .x1(x_05_037), .y0(x_06_036), .y1(x_06_037), .W(W009) );
    assign f_009 = x_06_036;
    assign f_041 = x_06_037;
    butt2 xx_05_010( .x0(x_05_020), .x1(x_05_021), .y0(x_06_020), .y1(x_06_021), .W(W010) );
    assign f_010 = x_06_020;
    assign f_042 = x_06_021;
    butt2 xx_05_011( .x0(x_05_052), .x1(x_05_053), .y0(x_06_052), .y1(x_06_053), .W(W011) );
    assign f_011 = x_06_052;
    assign f_043 = x_06_053;
    butt2 xx_05_012( .x0(x_05_012), .x1(x_05_013), .y0(x_06_012), .y1(x_06_013), .W(W012) );
    assign f_012 = x_06_012;
    assign f_044 = x_06_013;
    butt2 xx_05_013( .x0(x_05_044), .x1(x_05_045), .y0(x_06_044), .y1(x_06_045), .W(W013) );
    assign f_013 = x_06_044;
    assign f_045 = x_06_045;
    butt2 xx_05_014( .x0(x_05_028), .x1(x_05_029), .y0(x_06_028), .y1(x_06_029), .W(W014) );
    assign f_014 = x_06_028;
    assign f_046 = x_06_029;
    butt2 xx_05_015( .x0(x_05_060), .x1(x_05_061), .y0(x_06_060), .y1(x_06_061), .W(W015) );
    assign f_015 = x_06_060;
    assign f_047 = x_06_061;
    butt2 xx_05_016( .x0(x_05_002), .x1(x_05_003), .y0(x_06_002), .y1(x_06_003), .W(W016) );
    assign f_016 = x_06_002;
    assign f_048 = x_06_003;
    butt2 xx_05_017( .x0(x_05_034), .x1(x_05_035), .y0(x_06_034), .y1(x_06_035), .W(W017) );
    assign f_017 = x_06_034;
    assign f_049 = x_06_035;
    butt2 xx_05_018( .x0(x_05_018), .x1(x_05_019), .y0(x_06_018), .y1(x_06_019), .W(W018) );
    assign f_018 = x_06_018;
    assign f_050 = x_06_019;
    butt2 xx_05_019( .x0(x_05_050), .x1(x_05_051), .y0(x_06_050), .y1(x_06_051), .W(W019) );
    assign f_019 = x_06_050;
    assign f_051 = x_06_051;
    butt2 xx_05_020( .x0(x_05_010), .x1(x_05_011), .y0(x_06_010), .y1(x_06_011), .W(W020) );
    assign f_020 = x_06_010;
    assign f_052 = x_06_011;
    butt2 xx_05_021( .x0(x_05_042), .x1(x_05_043), .y0(x_06_042), .y1(x_06_043), .W(W021) );
    assign f_021 = x_06_042;
    assign f_053 = x_06_043;
    butt2 xx_05_022( .x0(x_05_026), .x1(x_05_027), .y0(x_06_026), .y1(x_06_027), .W(W022) );
    assign f_022 = x_06_026;
    assign f_054 = x_06_027;
    butt2 xx_05_023( .x0(x_05_058), .x1(x_05_059), .y0(x_06_058), .y1(x_06_059), .W(W023) );
    assign f_023 = x_06_058;
    assign f_055 = x_06_059;
    butt2 xx_05_024( .x0(x_05_006), .x1(x_05_007), .y0(x_06_006), .y1(x_06_007), .W(W024) );
    assign f_024 = x_06_006;
    assign f_056 = x_06_007;
    butt2 xx_05_025( .x0(x_05_038), .x1(x_05_039), .y0(x_06_038), .y1(x_06_039), .W(W025) );
    assign f_025 = x_06_038;
    assign f_057 = x_06_039;
    butt2 xx_05_026( .x0(x_05_022), .x1(x_05_023), .y0(x_06_022), .y1(x_06_023), .W(W026) );
    assign f_026 = x_06_022;
    assign f_058 = x_06_023;
    butt2 xx_05_027( .x0(x_05_054), .x1(x_05_055), .y0(x_06_054), .y1(x_06_055), .W(W027) );
    assign f_027 = x_06_054;
    assign f_059 = x_06_055;
    butt2 xx_05_028( .x0(x_05_014), .x1(x_05_015), .y0(x_06_014), .y1(x_06_015), .W(W028) );
    assign f_028 = x_06_014;
    assign f_060 = x_06_015;
    butt2 xx_05_029( .x0(x_05_046), .x1(x_05_047), .y0(x_06_046), .y1(x_06_047), .W(W029) );
    assign f_029 = x_06_046;
    assign f_061 = x_06_047;
    butt2 xx_05_030( .x0(x_05_030), .x1(x_05_031), .y0(x_06_030), .y1(x_06_031), .W(W030) );
    assign f_030 = x_06_030;
    assign f_062 = x_06_031;
    butt2 xx_05_031( .x0(x_05_062), .x1(x_05_063), .y0(x_06_062), .y1(x_06_063), .W(W031) );
    assign f_031 = x_06_062;
    assign f_063 = x_06_063;
endmodule
////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////
module butt2(y0,y1,x0,x1,W);
    input [31:0] x0,x1,W;
    output[31:0] y0,y1;

    wire [31:0] x11;

    assign x11 = mulc(x1, W);
    assign y0 = addc( x0, x11 );
    assign y1 = subc( x0, x11 );

    function [31:0] addc;
        input [31:0] a, b;
        reg [15:0] yr, yi;
        begin
            yr = a[31:16] + b[31:16];
            yi = a[15:0] + b[15:0];
            addc = {yr, yi};
        end
    endfunction
    function [31:0] subc;
        input [31:0] a, b;
        reg [15:0] yr, yi;
        begin
            yr = a[31:16] - b[31:16];
            yi = a[15:0] - b[15:0];
            subc = {yr, yi};
        end
    endfunction
    //  function [31:0] mulc;
    //    input [31:0] a, b;
    //    reg [15:0] yr, yi;
    //    begin
    //      yr = a[31:16]*b[31:16] - a[15:0]*b[15:0];
    //      yi = a[15:0]*b[31:16] + a[31:16]*b[15:0];
    //      mulc = {yr, yi};
    //    end
    //  endfunction
    function [31:0] mulc;
        input [31:0] a, b;
        reg [31:0] yr1, yr2, yi1, yi2;
        reg [15:0] ar, ai, br, bi, yyr1, yyr2, yyi1, yyi2, yr, yi;
        begin
            if( a[31] == 0 ) ar = a[31:16]; else ar = ~(a[31:16]-1);
            if( a[15] == 0 ) ai = a[15:0]; else ai = ~(a[15:0]-1);
            if( b[31] == 0 ) br = b[31:16]; else br = ~(b[31:16]-1);
            if( b[15] == 0 ) bi = b[15:0]; else bi = ~(b[15:0]-1);


            yr1 = ar * br;
            yr2 = ai * bi;

            yi1 = ar * bi;
            yi2 = ai * br;

            if( (a[31]^b[31])==0 ) yyr1 = yr1[26:11]; else yyr1 = ~yr1[26:11] + 1;
            if( (a[15]^b[15])==0 ) yyr2 = yr2[26:11]; else yyr2 = ~yr2[26:11] + 1;
            yr = yyr1 - yyr2;

            if( (a[31]^b[15])==0 ) yyi1 = yi1[26:11]; else yyi1 = ~yi1[26:11] + 1;
            if( (a[15]^b[31])==0 ) yyi2 = yi2[26:11]; else yyi2 = ~yi2[26:11] + 1;
            yi = yyi1 + yyi2;

            mulc = {yr, yi};
        end
    endfunction
endmodule
////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////
module top;
    wire [31:0]
                f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
                f_010,f_011,f_012,f_013,f_014,f_015,f_016,f_017,f_018,f_019,
                f_020,f_021,f_022,f_023,f_024,f_025,f_026,f_027,f_028,f_029,
                f_030,f_031,f_032,f_033,f_034,f_035,f_036,f_037,f_038,f_039,
                f_040,f_041,f_042,f_043,f_044,f_045,f_046,f_047,f_048,f_049,
                f_050,f_051,f_052,f_053,f_054,f_055,f_056,f_057,f_058,f_059,
                f_060,f_061,f_062,f_063;
    reg [31:0]
               x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
               x_010,x_011,x_012,x_013,x_014,x_015,x_016,x_017,x_018,x_019,
               x_020,x_021,x_022,x_023,x_024,x_025,x_026,x_027,x_028,x_029,
               x_030,x_031,x_032,x_033,x_034,x_035,x_036,x_037,x_038,x_039,
               x_040,x_041,x_042,x_043,x_044,x_045,x_046,x_047,x_048,x_049,
               x_050,x_051,x_052,x_053,x_054,x_055,x_056,x_057,x_058,x_059,
               x_060,x_061,x_062,x_063;
    reg [31:0]
               W000,W001,W002,W003,W004,W005,W006,W007,W008,W009,
               W010,W011,W012,W013,W014,W015,W016,W017,W018,W019,
               W020,W021,W022,W023,W024,W025,W026,W027,W028,W029,
               W030,W031;
    fft064 f(
             f_000,f_001,f_002,f_003,f_004,f_005,f_006,f_007,f_008,f_009,
             f_010,f_011,f_012,f_013,f_014,f_015,f_016,f_017,f_018,f_019,
             f_020,f_021,f_022,f_023,f_024,f_025,f_026,f_027,f_028,f_029,
             f_030,f_031,f_032,f_033,f_034,f_035,f_036,f_037,f_038,f_039,
             f_040,f_041,f_042,f_043,f_044,f_045,f_046,f_047,f_048,f_049,
             f_050,f_051,f_052,f_053,f_054,f_055,f_056,f_057,f_058,f_059,
             f_060,f_061,f_062,f_063,
             x_000,x_001,x_002,x_003,x_004,x_005,x_006,x_007,x_008,x_009,
             x_010,x_011,x_012,x_013,x_014,x_015,x_016,x_017,x_018,x_019,
             x_020,x_021,x_022,x_023,x_024,x_025,x_026,x_027,x_028,x_029,
             x_030,x_031,x_032,x_033,x_034,x_035,x_036,x_037,x_038,x_039,
             x_040,x_041,x_042,x_043,x_044,x_045,x_046,x_047,x_048,x_049,
             x_050,x_051,x_052,x_053,x_054,x_055,x_056,x_057,x_058,x_059,
             x_060,x_061,x_062,x_063,
             W000,W001,W002,W003,W004,W005,W006,W007,W008,W009,
             W010,W011,W012,W013,W014,W015,W016,W017,W018,W019,
             W020,W021,W022,W023,W024,W025,W026,W027,W028,W029,
             W030,W031);
    initial begin
        $dumpfile("fft.vcd");
        $dumpvars;
        W000 = { 16'b 0000100000000000, 16'b 0000000000000000 };
        W001 = { 16'b 0000011111110110, 16'b 1111111100111000 };
        W002 = { 16'b 0000011111011000, 16'b 1111111001110001 };
        W003 = { 16'b 0000011110100111, 16'b 1111110110101110 };
        W004 = { 16'b 0000011101100100, 16'b 1111110011110001 };
        W005 = { 16'b 0000011100001110, 16'b 1111110000111011 };
        W006 = { 16'b 0000011010100110, 16'b 1111101110001111 };
        W007 = { 16'b 0000011000101111, 16'b 1111101011101101 };
        W008 = { 16'b 0000010110101000, 16'b 1111101001011000 };
        W009 = { 16'b 0000010100010011, 16'b 1111100111010001 };
        W010 = { 16'b 0000010001110001, 16'b 1111100101011010 };
        W011 = { 16'b 0000001111000101, 16'b 1111100011110010 };
        W012 = { 16'b 0000001100001111, 16'b 1111100010011100 };
        W013 = { 16'b 0000001001010010, 16'b 1111100001011001 };
        W014 = { 16'b 0000000110001111, 16'b 1111100000101000 };
        W015 = { 16'b 0000000011001000, 16'b 1111100000001010 };
        W016 = { 16'b 0000000000000000, 16'b 1111100000000001 };
        W017 = { 16'b 1111111100111000, 16'b 1111100000001010 };
        W018 = { 16'b 1111111001110001, 16'b 1111100000101000 };
        W019 = { 16'b 1111110110101110, 16'b 1111100001011001 };
        W020 = { 16'b 1111110011110001, 16'b 1111100010011100 };
        W021 = { 16'b 1111110000111011, 16'b 1111100011110010 };
        W022 = { 16'b 1111101110001111, 16'b 1111100101011010 };
        W023 = { 16'b 1111101011101101, 16'b 1111100111010001 };
        W024 = { 16'b 1111101001011000, 16'b 1111101001011000 };
        W025 = { 16'b 1111100111010001, 16'b 1111101011101101 };
        W026 = { 16'b 1111100101011010, 16'b 1111101110001111 };
        W027 = { 16'b 1111100011110010, 16'b 1111110000111011 };
        W028 = { 16'b 1111100010011100, 16'b 1111110011110001 };
        W029 = { 16'b 1111100001011001, 16'b 1111110110101110 };
        W030 = { 16'b 1111100000101000, 16'b 1111111001110001 };
        W031 = { 16'b 1111100000001010, 16'b 1111111100111000 };
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_002 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_003 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_004 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_005 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_006 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_007 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_008 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_009 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_010 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_011 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_012 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_013 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_014 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_015 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_016 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_017 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_018 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_019 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_020 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_021 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_022 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_023 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_024 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_025 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_026 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_027 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_028 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_029 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_030 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_031 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_034 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_035 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_036 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_037 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_038 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_039 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_040 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_041 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_042 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_043 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_044 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_045 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_046 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_047 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_048 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_049 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_050 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_051 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_052 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_053 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_054 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_055 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_056 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_057 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_058 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_059 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_060 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_061 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_062 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_063 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_002 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_003 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_004 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_005 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_006 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_007 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_008 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_009 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_010 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_011 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_012 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_013 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_014 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_015 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_017 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_018 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_019 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_020 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_021 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_022 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_023 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_024 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_025 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_026 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_027 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_028 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_029 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_030 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_031 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_034 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_035 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_036 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_037 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_038 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_039 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_040 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_041 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_042 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_043 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_044 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_045 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_046 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_047 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_049 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_050 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_051 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_052 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_053 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_054 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_055 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_056 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_057 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_058 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_059 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_060 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_061 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_062 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_063 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_002 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_003 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_004 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_005 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_006 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_007 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_008 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_009 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_010 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_011 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_012 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_013 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_014 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_015 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_016 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_017 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_018 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_019 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_020 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_021 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_022 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_023 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_024 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_025 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_026 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_027 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_028 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_029 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_030 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_031 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_034 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_035 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_036 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_037 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_038 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_039 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_040 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_041 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_042 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_043 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_044 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_045 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_046 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_047 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_048 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_049 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_050 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_051 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_052 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_053 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_054 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_055 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_056 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_057 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_058 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_059 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_060 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_061 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_062 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_063 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_002 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_003 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_004 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_005 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_006 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_007 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_009 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_010 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_011 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_012 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_013 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_014 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_015 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_017 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_018 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_019 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_020 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_021 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_022 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_023 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_024 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_025 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_026 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_027 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_028 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_029 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_030 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_031 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_034 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_035 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_036 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_037 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_038 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_039 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_040 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_041 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_042 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_043 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_044 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_045 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_046 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_047 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_049 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_050 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_051 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_052 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_053 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_054 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_055 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_056 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_057 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_058 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_059 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_060 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_061 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_062 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_063 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_002 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_003 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_004 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_005 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_006 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_007 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_008 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_009 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_010 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_011 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_012 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_013 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_014 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_015 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_016 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_017 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_018 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_019 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_020 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_021 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_022 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_023 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_024 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_025 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_026 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_027 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_028 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_029 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_030 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_031 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_034 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_035 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_036 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_037 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_038 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_039 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_040 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_041 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_042 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_043 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_044 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_045 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_046 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_047 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_048 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_049 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_050 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_051 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_052 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_053 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_054 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_055 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_056 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_057 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_058 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_059 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_060 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_061 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_062 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_063 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_002 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_003 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_004 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_005 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_006 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_007 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_008 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_009 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_010 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_011 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_012 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_013 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_014 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_015 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_017 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_018 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_019 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_020 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_021 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_022 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_023 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_024 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_025 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_026 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_027 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_028 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_029 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_030 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_031 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_034 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_035 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_036 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_037 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_038 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_039 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_040 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_041 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_042 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_043 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_044 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_045 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_046 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_047 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_049 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_050 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_051 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_052 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_053 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_054 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_055 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_056 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_057 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_058 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_059 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_060 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_061 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_062 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_063 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_002 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_003 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_004 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_005 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_006 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_007 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_008 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_009 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_010 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_011 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_012 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_013 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_014 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_015 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_016 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_017 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_018 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_019 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_020 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_021 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_022 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_023 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_024 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_025 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_026 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_027 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_028 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_029 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_030 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_031 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_034 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_035 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_036 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_037 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_038 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_039 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_040 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_041 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_042 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_043 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_044 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_045 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_046 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_047 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_048 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_049 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_050 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_051 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_052 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_053 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_054 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_055 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_056 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_057 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_058 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_059 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_060 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_061 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_062 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_063 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_002 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_003 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_004 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_005 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_006 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_007 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_009 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_010 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_011 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_012 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_013 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_014 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_015 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_017 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_018 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_019 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_020 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_021 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_022 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_023 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_024 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_025 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_026 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_027 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_028 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_029 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_030 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_031 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_034 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_035 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_036 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_037 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_038 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_039 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_040 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_041 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_042 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_043 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_044 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_045 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_046 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_047 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_049 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_050 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_051 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_052 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_053 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_054 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_055 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_056 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_057 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_058 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_059 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_060 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_061 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_062 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_063 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_002 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_003 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_004 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_005 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_006 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_007 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_008 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_009 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_010 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_011 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_012 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_013 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_014 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_015 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_016 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_017 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_018 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_019 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_020 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_021 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_022 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_023 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_024 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_025 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_026 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_027 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_028 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_029 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_030 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_031 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_034 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_035 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_036 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_037 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_038 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_039 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_040 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_041 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_042 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_043 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_044 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_045 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_046 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_047 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_048 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_049 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_050 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_051 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_052 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_053 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_054 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_055 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_056 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_057 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_058 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_059 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_060 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_061 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_062 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_063 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_002 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_003 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_004 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_005 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_006 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_007 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_008 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_009 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_010 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_011 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_012 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_013 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_014 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_015 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_017 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_018 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_019 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_020 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_021 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_022 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_023 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_024 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_025 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_026 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_027 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_028 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_029 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_030 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_031 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_034 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_035 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_036 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_037 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_038 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_039 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_040 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_041 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_042 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_043 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_044 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_045 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_046 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_047 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_049 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_050 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_051 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_052 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_053 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_054 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_055 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_056 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_057 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_058 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_059 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_060 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_061 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_062 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_063 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_002 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_003 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_004 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_005 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_006 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_007 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_008 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_009 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_010 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_011 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_012 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_013 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_014 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_015 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_016 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_017 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_018 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_019 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_020 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_021 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_022 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_023 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_024 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_025 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_026 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_027 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_028 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_029 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_030 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_031 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_034 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_035 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_036 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_037 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_038 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_039 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_040 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_041 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_042 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_043 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_044 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_045 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_046 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_047 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_048 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_049 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_050 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_051 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_052 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_053 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_054 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_055 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_056 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_057 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_058 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_059 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_060 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_061 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_062 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_063 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_002 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_003 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_004 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_005 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_006 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_007 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_009 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_010 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_011 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_012 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_013 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_014 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_015 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_017 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_018 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_019 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_020 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_021 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_022 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_023 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_024 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_025 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_026 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_027 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_028 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_029 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_030 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_031 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_034 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_035 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_036 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_037 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_038 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_039 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_040 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_041 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_042 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_043 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_044 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_045 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_046 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_047 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_049 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_050 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_051 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_052 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_053 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_054 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_055 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_056 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_057 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_058 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_059 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_060 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_061 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_062 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_063 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_002 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_003 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_004 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_005 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_006 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_007 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_008 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_009 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_010 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_011 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_012 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_013 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_014 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_015 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_016 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_017 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_018 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_019 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_020 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_021 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_022 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_023 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_024 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_025 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_026 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_027 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_028 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_029 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_030 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_031 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_034 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_035 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_036 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_037 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_038 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_039 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_040 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_041 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_042 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_043 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_044 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_045 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_046 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_047 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_048 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_049 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_050 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_051 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_052 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_053 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_054 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_055 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_056 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_057 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_058 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_059 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_060 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_061 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_062 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_063 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_002 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_003 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_004 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_005 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_006 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_007 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_008 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_009 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_010 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_011 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_012 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_013 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_014 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_015 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_017 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_018 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_019 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_020 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_021 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_022 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_023 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_024 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_025 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_026 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_027 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_028 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_029 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_030 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_031 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_034 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_035 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_036 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_037 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_038 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_039 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_040 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_041 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_042 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_043 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_044 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_045 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_046 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_047 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_049 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_050 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_051 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_052 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_053 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_054 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_055 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_056 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_057 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_058 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_059 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_060 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_061 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_062 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_063 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_002 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_003 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_004 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_005 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_006 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_007 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_008 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_009 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_010 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_011 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_012 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_013 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_014 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_015 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_016 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_017 = { 16'b 1111111011111100, 16'b 0000000000000000 };   //  -0.127,  0.000
        x_018 = { 16'b 0000101000110011, 16'b 0000000000000000 };   //   1.275,  0.000
        x_019 = { 16'b 0000001100000100, 16'b 0000000000000000 };   //   0.377,  0.000
        x_020 = { 16'b 1111011001100101, 16'b 0000000000000000 };   //  -1.201,  0.000
        x_021 = { 16'b 1111101100011001, 16'b 0000000000000000 };   //  -0.613,  0.000
        x_022 = { 16'b 0000100010100101, 16'b 0000000000000000 };   //   1.081,  0.000
        x_023 = { 16'b 0000011010011001, 16'b 0000000000000000 };   //   0.825,  0.000
        x_024 = { 16'b 1111100010100110, 16'b 0000000000000000 };   //  -0.919,  0.000
        x_025 = { 16'b 1111011111110110, 16'b 0000000000000000 };   //  -1.005,  0.000
        x_026 = { 16'b 0000010111000111, 16'b 0000000000000000 };   //   0.722,  0.000
        x_027 = { 16'b 0000100100101100, 16'b 0000000000000000 };   //   1.146,  0.000
        x_028 = { 16'b 1111110000000110, 16'b 0000000000000000 };   //  -0.497,  0.000
        x_029 = { 16'b 1111011000001101, 16'b 0000000000000000 };   //  -1.244,  0.000
        x_030 = { 16'b 0000001000000111, 16'b 0000000000000000 };   //   0.254,  0.000
        x_031 = { 16'b 0000101001011001, 16'b 0000000000000000 };   //   1.294,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_033 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        x_034 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_035 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_036 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_037 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_038 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_039 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_040 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_041 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_042 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_043 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_044 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_045 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_046 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_047 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_048 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_049 = { 16'b 0000000100000100, 16'b 0000000000000000 };   //   0.127,  0.000
        x_050 = { 16'b 1111010111001101, 16'b 0000000000000000 };   //  -1.275,  0.000
        x_051 = { 16'b 1111110011111100, 16'b 0000000000000000 };   //  -0.377,  0.000
        x_052 = { 16'b 0000100110011011, 16'b 0000000000000000 };   //   1.201,  0.000
        x_053 = { 16'b 0000010011100111, 16'b 0000000000000000 };   //   0.613,  0.000
        x_054 = { 16'b 1111011101011011, 16'b 0000000000000000 };   //  -1.081,  0.000
        x_055 = { 16'b 1111100101100111, 16'b 0000000000000000 };   //  -0.825,  0.000
        x_056 = { 16'b 0000011101011010, 16'b 0000000000000000 };   //   0.919,  0.000
        x_057 = { 16'b 0000100000001010, 16'b 0000000000000000 };   //   1.005,  0.000
        x_058 = { 16'b 1111101000111001, 16'b 0000000000000000 };   //  -0.722,  0.000
        x_059 = { 16'b 1111011011010100, 16'b 0000000000000000 };   //  -1.146,  0.000
        x_060 = { 16'b 0000001111111010, 16'b 0000000000000000 };   //   0.497,  0.000
        x_061 = { 16'b 0000100111110011, 16'b 0000000000000000 };   //   1.244,  0.000
        x_062 = { 16'b 1111110111111001, 16'b 0000000000000000 };   //  -0.254,  0.000
        x_063 = { 16'b 1111010110100111, 16'b 0000000000000000 };   //  -1.294,  0.000
        #100
          $display( "f_000=%h", f_000);
        $display( "f_001=%h", f_001);
        $display( "f_002=%h", f_002);
        $display( "f_003=%h", f_003);
        $display( "f_004=%h", f_004);
        $display( "f_005=%h", f_005);
        $display( "f_006=%h", f_006);
        $display( "f_007=%h", f_007);
        $display( "f_008=%h", f_008);
        $display( "f_009=%h", f_009);
        $display( "f_010=%h", f_010);
        $display( "f_011=%h", f_011);
        $display( "f_012=%h", f_012);
        $display( "f_013=%h", f_013);
        $display( "f_014=%h", f_014);
        $display( "f_015=%h", f_015);
        $display( "f_016=%h", f_016);
        $display( "f_017=%h", f_017);
        $display( "f_018=%h", f_018);
        $display( "f_019=%h", f_019);
        $display( "f_020=%h", f_020);
        $display( "f_021=%h", f_021);
        $display( "f_022=%h", f_022);
        $display( "f_023=%h", f_023);
        $display( "f_024=%h", f_024);
        $display( "f_025=%h", f_025);
        $display( "f_026=%h", f_026);
        $display( "f_027=%h", f_027);
        $display( "f_028=%h", f_028);
        $display( "f_029=%h", f_029);
        $display( "f_030=%h", f_030);
        $display( "f_031=%h", f_031);
        $display( "f_032=%h", f_032);
        $display( "f_033=%h", f_033);
        $display( "f_034=%h", f_034);
        $display( "f_035=%h", f_035);
        $display( "f_036=%h", f_036);
        $display( "f_037=%h", f_037);
        $display( "f_038=%h", f_038);
        $display( "f_039=%h", f_039);
        $display( "f_040=%h", f_040);
        $display( "f_041=%h", f_041);
        $display( "f_042=%h", f_042);
        $display( "f_043=%h", f_043);
        $display( "f_044=%h", f_044);
        $display( "f_045=%h", f_045);
        $display( "f_046=%h", f_046);
        $display( "f_047=%h", f_047);
        $display( "f_048=%h", f_048);
        $display( "f_049=%h", f_049);
        $display( "f_050=%h", f_050);
        $display( "f_051=%h", f_051);
        $display( "f_052=%h", f_052);
        $display( "f_053=%h", f_053);
        $display( "f_054=%h", f_054);
        $display( "f_055=%h", f_055);
        $display( "f_056=%h", f_056);
        $display( "f_057=%h", f_057);
        $display( "f_058=%h", f_058);
        $display( "f_059=%h", f_059);
        $display( "f_060=%h", f_060);
        $display( "f_061=%h", f_061);
        $display( "f_062=%h", f_062);
        $display( "f_063=%h", f_063);
        x_000 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_001 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_002 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_003 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_004 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_005 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_006 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_007 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_008 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_009 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_010 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_011 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_012 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_013 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_014 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_015 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_016 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_017 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_018 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_019 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_020 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_021 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_022 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_023 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_024 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_025 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_026 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_027 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_028 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_029 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_030 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_031 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_032 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_033 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_034 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_035 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_036 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_037 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_038 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_039 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_040 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_041 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_042 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_043 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_044 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_045 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_046 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_047 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_048 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_049 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_050 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_051 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_052 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_053 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_054 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_055 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_056 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_057 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_058 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_059 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        x_060 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //  -0.000,  0.000
        x_061 = { 16'b 0000101001100110, 16'b 0000000000000000 };   //   1.300,  0.000
        x_062 = { 16'b 0000000000000000, 16'b 0000000000000000 };   //   0.000,  0.000
        x_063 = { 16'b 1111010110011010, 16'b 0000000000000000 };   //  -1.300,  0.000
        #100
          $finish;
    end
endmodule
