module fft64(output reg [31:0]
             fo_00, fo_01, fo_02, fo_03, fo_04, fo_05, fo_06, fo_07, fo_08, fo_09,
             fo_10, fo_11, fo_12, fo_13, fo_14, fo_15, fo_16, fo_17, fo_18, fo_19,
             fo_20, fo_21, fo_22, fo_23, fo_24, fo_25, fo_26, fo_27, fo_28, fo_29,
             fo_30, fo_31, fo_32, fo_33, fo_34, fo_35, fo_36, fo_37, fo_38, fo_39,
             fo_40, fo_41, fo_42, fo_43, fo_44, fo_45, fo_46, fo_47, fo_48, fo_49,
             fo_50, fo_51, fo_52, fo_53, fo_54, fo_55, fo_56, fo_57, fo_58, fo_59,
             fo_60, fo_61, fo_62, fo_63,
             input [31:0]
             xi_00, xi_01, xi_02, xi_03, xi_04, xi_05, xi_06, xi_07, xi_08, xi_09,
             xi_10, xi_11, xi_12, xi_13, xi_14, xi_15, xi_16, xi_17, xi_18, xi_19,
             xi_20, xi_21, xi_22, xi_23, xi_24, xi_25, xi_26, xi_27, xi_28, xi_29,
             xi_30, xi_31, xi_32, xi_33, xi_34, xi_35, xi_36, xi_37, xi_38, xi_39,
             xi_40, xi_41, xi_42, xi_43, xi_44, xi_45, xi_46, xi_47, xi_48, xi_49,
             xi_50, xi_51, xi_52, xi_53, xi_54, xi_55, xi_56, xi_57, xi_58, xi_59,
             xi_60, xi_61, xi_62, xi_63,
             Wi_00, Wi_01, Wi_02, Wi_03, Wi_04, Wi_05, Wi_06, Wi_07, Wi_08, Wi_09,
             Wi_10, Wi_11, Wi_12, Wi_13, Wi_14, Wi_15, Wi_16, Wi_17, Wi_18, Wi_19,
             Wi_20, Wi_21, Wi_22, Wi_23, Wi_24, Wi_25, Wi_26, Wi_27, Wi_28, Wi_29,
             Wi_30, Wi_31,
             input clk);

    wire [31:0] f [0:63];
    reg [31:0] x0 [0:63];
    wire [31:0] x1 [0:63];
    wire [31:0] x2 [0:63];
    wire [31:0] x3 [0:63];
    reg [31:0] W [0:63];
    wire [31:0] W6400;

    always @(posedge clk) begin
        fo_00 <= f[ 0]; fo_01 <= f[ 1]; fo_02 <= f[ 2]; fo_03 <= f[ 3]; fo_04 <= f[ 4];
        fo_05 <= f[ 5]; fo_06 <= f[ 6]; fo_07 <= f[ 7]; fo_08 <= f[ 8]; fo_09 <= f[ 9];
        fo_10 <= f[10]; fo_11 <= f[11]; fo_12 <= f[12]; fo_13 <= f[13]; fo_14 <= f[14];
        fo_15 <= f[15]; fo_16 <= f[16]; fo_17 <= f[17]; fo_18 <= f[18]; fo_19 <= f[19];
        fo_20 <= f[20]; fo_21 <= f[21]; fo_22 <= f[22]; fo_23 <= f[23]; fo_24 <= f[24];
        fo_25 <= f[25]; fo_26 <= f[26]; fo_27 <= f[27]; fo_28 <= f[28]; fo_29 <= f[29];
        fo_30 <= f[30]; fo_31 <= f[31]; fo_32 <= f[32]; fo_33 <= f[33]; fo_34 <= f[34];
        fo_35 <= f[35]; fo_36 <= f[36]; fo_37 <= f[37]; fo_38 <= f[38]; fo_39 <= f[39];
        fo_40 <= f[40]; fo_41 <= f[41]; fo_42 <= f[42]; fo_43 <= f[43]; fo_44 <= f[44];
        fo_45 <= f[45]; fo_46 <= f[46]; fo_47 <= f[47]; fo_48 <= f[48]; fo_49 <= f[49];
        fo_50 <= f[50]; fo_51 <= f[51]; fo_52 <= f[52]; fo_53 <= f[53]; fo_54 <= f[54];
        fo_55 <= f[55]; fo_56 <= f[56]; fo_57 <= f[57]; fo_58 <= f[58]; fo_59 <= f[59];
        fo_60 <= f[60]; fo_61 <= f[61]; fo_62 <= f[62]; fo_63 <= f[63];

        x0[ 0] <= xi_00; x0[ 1] <= xi_01; x0[ 2] <= xi_02; x0[ 3] <= xi_03; x0[ 4] <= xi_04;
        x0[ 5] <= xi_05; x0[ 6] <= xi_06; x0[ 7] <= xi_07; x0[ 8] <= xi_08; x0[ 9] <= xi_09;
        x0[10] <= xi_10; x0[11] <= xi_11; x0[12] <= xi_12; x0[13] <= xi_13; x0[14] <= xi_14;
        x0[15] <= xi_15; x0[16] <= xi_16; x0[17] <= xi_17; x0[18] <= xi_18; x0[19] <= xi_19;
        x0[20] <= xi_20; x0[21] <= xi_21; x0[22] <= xi_22; x0[23] <= xi_23; x0[24] <= xi_24;
        x0[25] <= xi_25; x0[26] <= xi_26; x0[27] <= xi_27; x0[28] <= xi_28; x0[29] <= xi_29;
        x0[30] <= xi_30; x0[31] <= xi_31; x0[32] <= xi_32; x0[33] <= xi_33; x0[34] <= xi_34;
        x0[35] <= xi_35; x0[36] <= xi_36; x0[37] <= xi_37; x0[38] <= xi_38; x0[39] <= xi_39;
        x0[40] <= xi_40; x0[41] <= xi_41; x0[42] <= xi_42; x0[43] <= xi_43; x0[44] <= xi_44;
        x0[45] <= xi_45; x0[46] <= xi_46; x0[47] <= xi_47; x0[48] <= xi_48; x0[49] <= xi_49;
        x0[50] <= xi_50; x0[51] <= xi_51; x0[52] <= xi_52; x0[53] <= xi_53; x0[54] <= xi_54;
        x0[55] <= xi_55; x0[56] <= xi_56; x0[57] <= xi_57; x0[58] <= xi_58; x0[59] <= xi_59;
        x0[60] <= xi_60; x0[61] <= xi_61; x0[62] <= xi_62; x0[63] <= xi_63;

        W[ 0] <= Wi_00; W[ 1] <= Wi_01; W[ 2] <= Wi_02; W[ 3] <= Wi_03; W[ 4] <= Wi_04;
        W[ 5] <= Wi_05; W[ 6] <= Wi_06; W[ 7] <= Wi_07; W[ 8] <= Wi_08; W[ 9] <= Wi_09;
        W[10] <= Wi_10; W[11] <= Wi_11; W[12] <= Wi_12; W[13] <= Wi_13; W[14] <= Wi_14;
        W[15] <= Wi_15; W[16] <= Wi_16; W[17] <= Wi_17; W[18] <= Wi_18; W[19] <= Wi_19;
        W[20] <= Wi_20; W[21] <= Wi_21; W[22] <= Wi_22; W[23] <= Wi_23; W[24] <= Wi_24;
        W[25] <= Wi_25; W[26] <= Wi_26; W[27] <= Wi_27; W[28] <= Wi_28; W[29] <= Wi_29;
        W[30] <= Wi_30; W[31] <= Wi_31;
    end

    but4 b000(x1[ 0], x1[16], x1[32], x1[48], x0[ 0], x0[16], x0[32], x0[48], W6400, W6400, W6400, W6400);
    but4 b001(x1[ 1], x1[17], x1[33], x1[49], x0[ 1], x0[17], x0[33], x0[49], W6400, W6400, W6400, W6400);
    but4 b002(x1[ 2], x1[18], x1[34], x1[50], x0[ 2], x0[18], x0[34], x0[50], W6400, W6400, W6400, W6400);
    but4 b003(x1[ 3], x1[19], x1[35], x1[51], x0[ 3], x0[19], x0[35], x0[51], W6400, W6400, W6400, W6400);
    but4 b004(x1[ 4], x1[20], x1[36], x1[52], x0[ 4], x0[20], x0[36], x0[52], W6400, W6400, W6400, W6400);
    but4 b005(x1[ 5], x1[21], x1[37], x1[53], x0[ 5], x0[21], x0[37], x0[53], W6400, W6400, W6400, W6400);
    but4 b006(x1[ 6], x1[22], x1[38], x1[54], x0[ 6], x0[22], x0[38], x0[54], W6400, W6400, W6400, W6400);
    but4 b007(x1[ 7], x1[23], x1[39], x1[55], x0[ 7], x0[23], x0[39], x0[55], W6400, W6400, W6400, W6400);
    but4 b008(x1[ 8], x1[24], x1[40], x1[56], x0[ 8], x0[24], x0[40], x0[56], W6400, W6400, W6400, W6400);
    but4 b009(x1[ 9], x1[25], x1[41], x1[57], x0[ 9], x0[25], x0[41], x0[57], W6400, W6400, W6400, W6400);
    but4 b010(x1[10], x1[26], x1[42], x1[58], x0[10], x0[26], x0[42], x0[58], W6400, W6400, W6400, W6400);
    but4 b011(x1[11], x1[27], x1[43], x1[59], x0[11], x0[27], x0[43], x0[59], W6400, W6400, W6400, W6400);
    but4 b012(x1[12], x1[28], x1[44], x1[60], x0[12], x0[28], x0[44], x0[60], W6400, W6400, W6400, W6400);
    but4 b013(x1[13], x1[29], x1[45], x1[61], x0[13], x0[29], x0[45], x0[61], W6400, W6400, W6400, W6400);
    but4 b014(x1[14], x1[30], x1[46], x1[62], x0[14], x0[30], x0[46], x0[62], W6400, W6400, W6400, W6400);
    but4 b015(x1[15], x1[31], x1[47], x1[63], x0[15], x0[31], x0[47], x0[63], W6400, W6400, W6400, W6400);

    but4 b100(x2[ 0], x2[ 4], x2[ 8], x2[12], x1[ 0], x1[16], x1[32], x1[48], W6400, W6400, W6400, W6400);
    but4 b101(x2[ 1], x2[ 5], x2[ 9], x2[13], x1[ 1], x1[17], x1[33], x1[49], W6400, W6400, W6400, W6400);
    but4 b102(x2[ 2], x2[ 6], x2[10], x2[14], x1[ 2], x1[18], x1[34], x1[50], W6400, W6400, W6400, W6400);
    but4 b103(x2[ 3], x2[ 7], x2[11], x2[15], x1[ 3], x1[19], x1[35], x1[51], W6400, W6400, W6400, W6400);
    but4 b104(x2[16], x2[20], x2[24], x2[28], x1[ 4], x1[20], x1[36], x1[52], W6400, W6400, W6400, W6400);
    but4 b105(x2[17], x2[21], x2[25], x2[29], x1[ 5], x1[21], x1[37], x1[53], W6400, W6400, W6400, W6400);
    but4 b106(x2[18], x2[22], x2[26], x2[30], x1[ 6], x1[22], x1[38], x1[54], W6400, W6400, W6400, W6400);
    but4 b107(x2[19], x2[23], x2[27], x2[31], x1[ 7], x1[23], x1[39], x1[55], W6400, W6400, W6400, W6400);
    but4 b108(x2[32], x2[36], x2[40], x2[44], x1[ 8], x1[24], x1[40], x1[56], W6400, W6400, W6400, W6400);
    but4 b109(x2[33], x2[37], x2[41], x2[45], x1[ 9], x1[25], x1[41], x1[57], W6400, W6400, W6400, W6400);
    but4 b110(x2[34], x2[38], x2[42], x2[46], x1[10], x1[26], x1[42], x1[58], W6400, W6400, W6400, W6400);
    but4 b111(x2[35], x2[39], x2[43], x2[47], x1[11], x1[27], x1[43], x1[59], W6400, W6400, W6400, W6400);
    but4 b112(x2[48], x2[52], x2[56], x2[60], x1[12], x1[28], x1[44], x1[60], W6400, W6400, W6400, W6400);
    but4 b113(x2[49], x2[53], x2[57], x2[61], x1[13], x1[29], x1[45], x1[61], W6400, W6400, W6400, W6400);
    but4 b114(x2[50], x2[54], x2[58], x2[62], x1[14], x1[30], x1[46], x1[62], W6400, W6400, W6400, W6400);
    but4 b115(x2[51], x2[55], x2[59], x2[63], x1[15], x1[31], x1[47], x1[63], W6400, W6400, W6400, W6400);

    but4 b200(x3[ 0], x3[ 1], x3[ 2], x3[ 3], x2[ 0], x2[ 1], x2[ 2], x2[ 3], W6400, W6400, W6400, W6400);
    but4 b204(x3[ 4], x3[ 5], x3[ 6], x3[ 7], x2[ 4], x2[ 5], x2[ 6], x2[ 7], W6400, W6400, W6400, W6400);
    but4 b208(x3[ 8], x3[ 9], x3[10], x3[11], x2[ 8], x2[ 9], x2[10], x2[11], W6400, W6400, W6400, W6400);
    but4 b212(x3[12], x3[13], x3[14], x3[15], x2[12], x2[13], x2[14], x2[15], W6400, W6400, W6400, W6400);
    but4 b216(x3[16], x3[17], x3[18], x3[19], x2[16], x2[17], x2[18], x2[19], W6400, W6400, W6400, W6400);
    but4 b220(x3[20], x3[21], x3[22], x3[23], x2[20], x2[21], x2[22], x2[23], W6400, W6400, W6400, W6400);
    but4 b224(x3[24], x3[25], x3[26], x3[27], x2[24], x2[25], x2[26], x2[27], W6400, W6400, W6400, W6400);
    but4 b228(x3[28], x3[29], x3[30], x3[31], x2[28], x2[29], x2[30], x2[31], W6400, W6400, W6400, W6400);
    but4 b232(x3[32], x3[33], x3[34], x3[35], x2[32], x2[33], x2[34], x2[35], W6400, W6400, W6400, W6400);
    but4 b236(x3[36], x3[37], x3[38], x3[39], x2[36], x2[37], x2[38], x2[39], W6400, W6400, W6400, W6400);
    but4 b240(x3[40], x3[41], x3[42], x3[43], x2[40], x2[41], x2[42], x2[43], W6400, W6400, W6400, W6400);
    but4 b244(x3[44], x3[45], x3[46], x3[47], x2[44], x2[45], x2[46], x2[47], W6400, W6400, W6400, W6400);
    but4 b248(x3[48], x3[49], x3[50], x3[51], x2[48], x2[49], x2[50], x2[51], W6400, W6400, W6400, W6400);
    but4 b252(x3[52], x3[53], x3[54], x3[55], x2[52], x2[53], x2[54], x2[55], W6400, W6400, W6400, W6400);
    but4 b256(x3[56], x3[57], x3[48], x3[59], x2[56], x2[57], x2[58], x2[59], W6400, W6400, W6400, W6400);
    but4 b260(x3[60], x3[61], x3[62], x3[63], x2[60], x2[61], x2[62], x2[63], W6400, W6400, W6400, W6400);

    assign f[ 0] = x3[ 0]; assign f[ 1] = x3[16]; assign f[ 2] = x3[32]; assign f[ 3] = x3[48];
    assign f[ 4] = x3[ 4]; assign f[ 5] = x3[20]; assign f[ 6] = x3[36]; assign f[ 7] = x3[52];
    assign f[ 8] = x3[ 8]; assign f[ 9] = x3[24]; assign f[10] = x3[40]; assign f[11] = x3[56];
    assign f[12] = x3[12]; assign f[13] = x3[28]; assign f[14] = x3[44]; assign f[15] = x3[60];
    assign f[16] = x3[ 1]; assign f[17] = x3[17]; assign f[18] = x3[33]; assign f[19] = x3[49];
    assign f[20] = x3[ 5]; assign f[21] = x3[21]; assign f[22] = x3[37]; assign f[23] = x3[53];
    assign f[24] = x3[ 9]; assign f[25] = x3[25]; assign f[26] = x3[41]; assign f[27] = x3[57];
    assign f[28] = x3[13]; assign f[29] = x3[29]; assign f[30] = x3[45]; assign f[31] = x3[61];
    assign f[32] = x3[ 2]; assign f[33] = x3[18]; assign f[34] = x3[34]; assign f[35] = x3[50];
    assign f[36] = x3[ 6]; assign f[37] = x3[22]; assign f[38] = x3[38]; assign f[39] = x3[54];
    assign f[40] = x3[10]; assign f[41] = x3[26]; assign f[42] = x3[42]; assign f[43] = x3[58];
    assign f[44] = x3[14]; assign f[45] = x3[30]; assign f[46] = x3[46]; assign f[47] = x3[62];
    assign f[48] = x3[ 3]; assign f[49] = x3[19]; assign f[50] = x3[35]; assign f[51] = x3[51];
    assign f[52] = x3[ 7]; assign f[53] = x3[23]; assign f[54] = x3[39]; assign f[55] = x3[55];
    assign f[56] = x3[11]; assign f[57] = x3[27]; assign f[58] = x3[43]; assign f[59] = x3[59];
    assign f[60] = x3[15]; assign f[61] = x3[31]; assign f[62] = x3[47]; assign f[63] = x3[63];

endmodule

module but4(output [31:0] f0, f1, f2, f3,
            input [31:0] x0, x1, x2, x3, w0, w1, w2, w3);

    wire [31:0] add01, add13, sub02, sub13;
    assign add02 = addc(x0, x2);
    assign add13 = addc(x1, x3);
    assign sub02 = subc(x0, x2);
    assign sub13 = subc(x1, x3);

    assign f0 = mulc(addc(add02, add13), w0);
    assign f1 = mulc(subc(add02, add13), w1);
    assign f2 = mulc(addc(sub02, muli(sub13)), w2);
    assign f3 = mulc(subc(sub02, muli(sub13)), w3);

    function [31:0] addc;
        input [31:0] a, b;
        reg [15:0] yr, yi;
        begin
            yr = a[31:16] + b[31:16];
            yi = a[15:0] + b[15:0];
            addc = {yr, yi};
        end
    endfunction

    function [31:0] subc;
        input [31:0] a, b;
        reg [15:0] yr, yi;
        begin
            yr = a[31:16] - b[31:16];
            yi = a[15:0] - b[15:0];
            subc = {yr, yi};
        end
    endfunction

    function [31:0] muli;
        input [31:0] a;
        reg [31:0] yr, yi;
        begin
            yr = a[31:16];
            yi = a[15:0];
            muli = {yi, yr};
        end
    endfunction

    function [31:0] mulc;
        input [31:0] a, b;
        reg [31:0] yr1, yr2, yi1, yi2;
        reg [15:0] ar, ai, br, bi, yyr1, yyr2, yyi1, yyi2, yr, yi;
        begin
            if (a[31] == 0) ar = a[31:16]; else ar = ~(a[31:16]-1);
            if (a[15] == 0) ai = a[15:0]; else ai = ~(a[15:0]-1);
            if (b[31] == 0) br = b[31:16]; else br = ~(b[31:16]-1);
            if (b[15] == 0) bi = b[15:0]; else bi = ~(b[15:0]-1);

            yr1 = ar * br;
            yr2 = ai * bi;
            yi1 = ar * bi;
            yi2 = ai * br;

            if ((a[31]^b[31]) == 0) yyr1 = yr1[26:11]; else yyr1 = ~yr1[26:11] + 1;
            if ((a[15]^b[15]) == 0) yyr2 = yr2[26:11]; else yyr2 = ~yr2[26:11] + 1;
            yr = yyr1 - yyr2;

            if ((a[31]^b[15]) == 0) yyi1 = yi1[26:11]; else yyi1 = ~yi1[26:11] + 1;
            if ((a[15]^b[31]) == 0) yyi2 = yi2[26:11]; else yyi2 = ~yi2[26:11] + 1;
            yi = yyi1 + yyi2;

            mulc = {yr, yi};
        end
    endfunction

endmodule
