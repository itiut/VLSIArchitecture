module processor(input clk,
                 input n_rst);
endmodule
